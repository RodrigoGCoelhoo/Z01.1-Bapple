--
-- Elementos de Sistemas - Aula 5 - Logica Combinacional
-- Rafael . Corsi @ insper . edu . br
--
-- Arquivo exemplo para acionar os LEDs e ler os bottoes
-- da placa DE0-CV utilizada no curso de elementos de
-- sistemas do 3s da eng. da computacao

----------------------------
-- Bibliotecas ieee       --
----------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

----------------------------
-- Entrada e saidas do bloco
----------------------------
entity TopLevel is
	port(
		CLOCK_50 : in  std_logic;
		SW       : in  std_logic_vector(9 downto 0);
		signal x	: buffer std_logic;
		signal y	: buffer std_logic;
		signal z	: buffer std_logic;
		a 			: out std_logic;
		LEDR     : out std_logic_vector(9 downto 0)
		
	);
end entity;

----------------------------
-- Implementacao do bloco --
----------------------------
architecture rtl of TopLevel is

--------------
-- signals
--------------
	
---------------
-- implementacao
---------------
begin

	x <= SW(0);
	y <= SW(1);
	z <= SW(2);
	
	a <= ((not((x and y) or y)) or (not(x and y and z)));
	
	
	
		
	

end rtl;
